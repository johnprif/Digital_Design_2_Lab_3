library verilog;
use verilog.vl_types.all;
entity AccumulatorLCD_vlg_vec_tst is
end AccumulatorLCD_vlg_vec_tst;
