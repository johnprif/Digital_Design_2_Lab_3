library verilog;
use verilog.vl_types.all;
entity Fibonacci_vlg_vec_tst is
end Fibonacci_vlg_vec_tst;
