library verilog;
use verilog.vl_types.all;
entity my_register_vlg_vec_tst is
end my_register_vlg_vec_tst;
